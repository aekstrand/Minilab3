module tb_spart(
    input clk,
    input rst_n,
    input rxd,
    input [7:0] rdata,
    output txd,
    output [7:0] tdata
);

endmodule