module tb_spart(
    input clk,
    input rst_n,
    input rxd,
    output [7:0] rdata,
    output txd,
    input [7:0] tdata,
    input rx_done,
    input start_transmission
);

endmodule